pBAV       �j ��   @  �����F?   ���������F?   ���������F?   ���������F?   ���������F?   ���������F?   ���������F?   ���������F?   ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������  �F    ��������
 @H        �����_   � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � � 
 @H        �����  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � 
 @H        �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � 
 @H        �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � 
 @H        �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � 
 @H        �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � 
 @H        �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � 
 @H        �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �   ���	FL(�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              