pBAV        � ��   @  ����d��@�  ��������d��@�  ��������d��@�  ��������d��@�  ��������d��@�  ��������d��@�  ��������d��@�  ��������d��@�  ��������d��@�  ��������d��@�  ��������d��@�  ��������d��@�  ����������@�  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  D( ((      �����_   � � � �   @$ $$      �����_   � � � �  2* **      �����_   � � � �  H311      �����_   � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �  @T  x      �����_  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  @`  x      �����_  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �   @<  x      �����_  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �   @<  x      �����_  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  @T x      �����_  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  @` x      �����_  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  @K  x      �����_ 	 � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  @H  x      �����_ 
 � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �   @H  x      �����	  � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �   @<  x      �����_
  � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �   @<  x      �����_  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  @T  x      �����_  � � � �  @T  x      �����_  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �   �T��X����F  �j	�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  