pBAV       � ��   @  ������?   ����������?   ����������?   ����������?   ����������?   ����������?   ����������?   ����������?   ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������
 @H        �����_   � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � � 
 @H        �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � 
 @H        �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � 
 @H        �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � 
 @H        �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � 
 @H        �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � 
 @H        �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � 
 @H        �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �   R�	|
22�Z�	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              