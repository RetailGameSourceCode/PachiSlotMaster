pBAV       Ў ��   @  ������?   ����������?   ����������?   ����������?   ����������?   ����������?   ����������?   ����������?   ����������?   ����������?   ����������?   ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������
 @H        �����_   � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � � 
 @H        �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � 
 @H        �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � 
 @H        �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � 
 @H        �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � 
 @H        �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � 
 @H        �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � 
 @H        �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � 
 @<        �����_ 	 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � 
 @H        �����_	 
 � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � � 
 @T        �����_
  � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �   �2X � �	�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        